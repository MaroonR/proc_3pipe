`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:22:55 04/27/2015 
// Design Name: 
// Module Name:    instruction_fetch 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: loads the instruction from memory, increments the program counter
// 				 by four, feeds into ld_st reg at the end
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module instruction_fetch(
    );

	HW8_n_bit_PC PC()
	//hw1_BFA_gate ADD4(a, b, cin, s, cout) not even sure we need this
endmodule
